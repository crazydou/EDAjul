LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY KEYBOARD_EV IS
PORT(
  CLK  : IN  STD_LOGIC;
    V  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);--SUPPORTING THAT THERE IS ONLY ONE SIGNAL
    O  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);--GIVE THE TRANSFORMATION OF THE MATRIX KEYBOARD IN BINARY
	D  : OUT STD_LOGIC;--INFORM THE STATE 
    H  : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)--TO SCAN THE KEYBOARD
    );
END ENTITY KEYBOARD_EV;
ARCHITECTURE BEHAVR OF KEYBOARD_EV IS
TYPE STATE_TYPE IS (S1,S2,S3,S4);
SIGNAL STATE:STATE_TYPE;
BEGIN
P1: PROCESS(CLK,V)
BEGIN
IF V=0 THEN
   IF (CLK'EVENT AND CLK='1') THEN
          CASE STATE IS
          WHEN S1=> STATE<=S2;
          WHEN S2=> STATE<=S3;
          WHEN S3=> STATE<=S4;  
          WHEN S4=> STATE<=S1; 
          END CASE;
   END IF;
END IF;
END PROCESS;
P2: PROCESS(STATE)
BEGIN
CASE STATE IS
WHEN S1=> H<="1000";
WHEN S2=> H<="0100";
WHEN S3=> H<="0010";  
WHEN S4=> H<="0001"; 
END CASE;
END PROCESS;
P3: PROCESS(V)
VARIABLE P : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
IF V>0 THEN
   IF V="1000" THEN
      CASE STATE IS
      WHEN S1=> P :="0001";D<='1';
      WHEN S2=> P :="0010";D<='1';
      WHEN S3=> P :="0011";D<='1';
      WHEN S4=> P :="0100";D<='1';
      END CASE;
   ELSIF V="0100" THEN
      CASE STATE IS
      WHEN S1=> P :="0101";D<='1';
      WHEN S2=> P :="0110";D<='1';
      WHEN S3=> P :="0111";D<='1';
      WHEN S4=> P :="1000";D<='1';
      END CASE;
   ELSIF V="0010" THEN
      CASE STATE IS
      WHEN S1=> P :="1001";D<='1';
      WHEN S2=> P :="1010";D<='1';
      WHEN S3=> P :="1011";D<='1';
      WHEN S4=> P :="1100";D<='1';
	  END CASE;
   ELSIF V="0001" THEN
	  CASE STATE IS
	  WHEN S1=> P :="0000";D<='1';
	  WHEN S2=> P :="1101";D<='1';
	  WHEN S3=> P :="1110";D<='1';
	  WHEN S4=> P :="0000";D<='0';
	  END CASE; 
   END IF;
   ELSE P:="0000";D<='0';
END IF;
O<=P;
END PROCESS;
END BEHAVR;
