--THE KEYBOARDSCAN VHDL FILE--
--By Wang Qin 
--2013/5/20 1:26
--AllCapClass STYLE
--END 

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY KEYSCAN IS                                  --ENTITY for KEYSCAN
	PORT(
		CLK:IN STD_LOGIC;				
		KBCOL:IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		KBROW:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		KBDOWN:OUT STD_LOGIC;
		KBDATA:OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END KEYSCAN;

ARCHITECTURE ONE OF KEYSCAN IS
SIGNAL CLK_NEW:STD_LOGIC;
SIGNAL ROWREG:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CON:STD_LOGIC_VECTOR(7 DOWNTO 0);

COMPONENT clkdiv is
--  generic(N: integer:=10);         					--N is the slip rate  /copied from clkdiv.vhd/          
  port(
        clkin: IN std_logic;
        clkout: OUT std_logic
        );
END COMPONENT;

BEGIN
U1: clkdiv PORT MAP(clkin=>CLK,clkout=>CLK_NEW);       	--slip the clock

U2:PROCESS(CLK_NEW)										--generate the rowscan signal
	BEGIN
	IF CLK_NEW'EVENT AND CLK_NEW='1' THEN
		CASE ROWREG IS 
			WHEN "0001"=>ROWREG<="0010";
			WHEN "0010"=>ROWREG<="0100";
			WHEN "0100"=>ROWREG<="1000";
			WHEN "1000"=>ROWREG<="0001";
			WHEN OTHERS=>ROWREG<="0001";
		END CASE;
	END IF;
END PROCESS U2;

KBROW<=ROWREG;
CON<=ROWREG&KBCOL;

U3:PROCESS(CLK_NEW,CON)
	BEGIN
	IF CLK_NEW'EVENT AND CLK_NEW='1' THEN
		CASE CON IS 
			WHEN "00010001"=>
			KBDATA<="0001";
			KBDOWN<='1';
			WHEN "00100001"=>
			KBDATA<="0010";
			KBDOWN<='1';
			WHEN "01000001"=>
			KBDATA<="0011";
			KBDOWN<='1';
			WHEN "10000001"=>
			KBDATA<="0100";
			KBDOWN<='1';
			WHEN "00010010"=>
			KBDATA<="0101";
			KBDOWN<='1';
			WHEN "00100010"=>
			KBDATA<="0110";
			KBDOWN<='1';
			WHEN "01000010"=>
			KBDATA<="0111";
			KBDOWN<='1';
			WHEN "10000010"=>
			KBDATA<="1000";
			KBDOWN<='1';
			WHEN "00010100"=>
			KBDATA<="1001";
			KBDOWN<='1';
			WHEN "00011000"=>
			KBDATA<="0000";
			KBDOWN<='1';
			WHEN "00100100"=>
			KBDATA<="1010";
			KBDOWN<='1';
			WHEN "01000100"=>
			KBDATA<="1011";
			KBDOWN<='1';
			WHEN "10000100"=>
			KBDATA<="1100";
			KBDOWN<='1';
			WHEN "00101000"=>
			KBDATA<="1101";
			KBDOWN<='1';
			WHEN "01001000"=>
			KBDATA<="1110";
			KBDOWN<='1';
			WHEN "10001000"=>
			KBDATA<="1111";
			KBDOWN<='1';
		WHEN OTHERS=>KBDOWN<='0';
		END CASE;
	END IF;
	END PROCESS;
END ONE;
